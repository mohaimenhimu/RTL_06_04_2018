`define TX